-------------------------------------------------------------------------
-- Justin Sebahar
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------
-- decoder5t32
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 5-to-32 decoder implemented with dataflow

-- 9/4/24
-------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ENTITY decoder5t32 IS
	PORT (
		i_IN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		i_EN : IN STD_LOGIC;
		o_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END decoder5t32;

ARCHITECTURE dataflow OF decoder5t32 IS
BEGIN
	o_OUT <= "00000000000000000000000000000000" WHEN (i_EN = '0') ELSE
		"00000000000000000000000000000001" WHEN (i_IN = "00000") ELSE
		"00000000000000000000000000000010" WHEN (i_IN = "00001") ELSE
		"00000000000000000000000000000100" WHEN (i_IN = "00010") ELSE
		"00000000000000000000000000001000" WHEN (i_IN = "00011") ELSE
		"00000000000000000000000000010000" WHEN (i_IN = "00100") ELSE
		"00000000000000000000000000100000" WHEN (i_IN = "00101") ELSE
		"00000000000000000000000001000000" WHEN (i_IN = "00110") ELSE
		"00000000000000000000000010000000" WHEN (i_IN = "00111") ELSE
		"00000000000000000000000100000000" WHEN (i_IN = "01000") ELSE
		"00000000000000000000001000000000" WHEN (i_IN = "01001") ELSE
		"00000000000000000000010000000000" WHEN (i_IN = "01010") ELSE
		"00000000000000000000100000000000" WHEN (i_IN = "01011") ELSE
		"00000000000000000001000000000000" WHEN (i_IN = "01100") ELSE
		"00000000000000000010000000000000" WHEN (i_IN = "01101") ELSE
		"00000000000000000100000000000000" WHEN (i_IN = "01110") ELSE
		"00000000000000001000000000000000" WHEN (i_IN = "01111") ELSE
		"00000000000000010000000000000000" WHEN (i_IN = "10000") ELSE
		"00000000000000100000000000000000" WHEN (i_IN = "10001") ELSE
		"00000000000001000000000000000000" WHEN (i_IN = "10010") ELSE
		"00000000000010000000000000000000" WHEN (i_IN = "10011") ELSE
		"00000000000100000000000000000000" WHEN (i_IN = "10100") ELSE
		"00000000001000000000000000000000" WHEN (i_IN = "10101") ELSE
		"00000000010000000000000000000000" WHEN (i_IN = "10110") ELSE
		"00000000100000000000000000000000" WHEN (i_IN = "10111") ELSE
		"00000001000000000000000000000000" WHEN (i_IN = "11000") ELSE
		"00000010000000000000000000000000" WHEN (i_IN = "11001") ELSE
		"00000100000000000000000000000000" WHEN (i_IN = "11010") ELSE
		"00001000000000000000000000000000" WHEN (i_IN = "11011") ELSE
		"00010000000000000000000000000000" WHEN (i_IN = "11100") ELSE
		"00100000000000000000000000000000" WHEN (i_IN = "11101") ELSE
		"01000000000000000000000000000000" WHEN (i_IN = "11110") ELSE
		"10000000000000000000000000000000" WHEN (i_IN = "11111") ELSE
		"00000000000000000000000000000000";

END dataflow;